library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.STD_LOGIC_UNSIGNED.all;
use IEEE.STD_LOGIC_ARITH.all;


entity AFISARE is
	port(ETAJ:in STD_LOGIC_VECTOR(3 downto 0);
	CLOCK:in STD_LOGIC;
	CATOD:out STD_LOGIC_VECTOR(6 downto 0);
	ANOD:out STD_LOGIC_VECTOR(3 downto 0));
end entity AFISARE;

architecture F_AFISARE of AFISARE is
signal CIFRA_ZECI,CIFRA_UNITATI:STD_LOGIC_VECTOR(3 downto 0);
signal CLOCK_DIVIZAT:STD_LOGIC;

begin
	A1:entity work.DECODIFICATOR(F_DECODIFICATOR) PORT MAP (ETAJ,CIFRA_ZECI,CIFRA_UNITATI);
	A2:entity work.AFISOR(F_AFISOR) PORT MAP (CLOCK,"1111",CIFRA_ZECI,CIFRA_UNITATI,"1111",ANOD,CATOD);
end architecture F_AFISARE;	



	
