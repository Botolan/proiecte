library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.STD_LOGIC_UNSIGNED.all;
--use IEEE.STD_LOGIC_ARITH.all;
use ieee.numeric_std.all;



entity OPRIRE is
	port(ETAJ_CURENT,ETAJ_MINIM_MAXIM:in STD_LOGIC_VECTOR(3 downto 0);
	INFORMATIE_IN:in STD_LOGIC_VECTOR(1 downto 0);
	SENS,CLOCK,SENZOR_USA,SENZOR_GREUTATE:in STD_LOGIC;
	ENABLE_NUMARATOR_OUT,ENABLE_DELETE:out STD_LOGIC);	
end entity OPRIRE;


architecture F_OPRIRE of OPRIRE is

signal REZULTATE_VALIDARE:STD_LOGIC_VECTOR(1 downto 0) := "11";
signal ENABLE_NUMARATOR,DELETE,CLOCK_DIVIZAT:STD_LOGIC := '0';


begin
	
	V1:entity work.VALIDARE(F_VALIDARE) PORT MAP (ETAJ_CURENT,ETAJ_MINIM_MAXIM,INFORMATIE_IN,SENS,CLOCK,DELETE,REZULTATE_VALIDARE);
	V2:entity work.TIMER_USA(F_TIMER_USA) PORT MAP (REZULTATE_VALIDARE,ETAJ_MINIM_MAXIM,CLOCK_DIVIZAT,SENZOR_USA,SENZOR_GREUTATE,ENABLE_NUMARATOR);
	V3:entity work.DIVIZOR_1_SEC(F_DIVIZOR_1_SEC) PORT MAP (CLOCK,CLOCK_DIVIZAT);
	
	
	ENABLE_NUMARATOR_OUT <= 
	'1' when REZULTATE_VALIDARE /= "01" and REZULTATE_VALIDARE /= "10" and ENABLE_NUMARATOR = '1' and ETAJ_MINIM_MAXIM /= "1111" else
	'0';
	
	ENABLE_DELETE <= DELETE and not(ENABLE_NUMARATOR);
	
	 
	
end architecture F_OPRIRE;



