library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.STD_LOGIC_UNSIGNED.all;
--use IEEE.STD_LOGIC_ARITH.all;
use ieee.numeric_std.all;


entity AUTOMAT is
	port(INFORMATIE_IN:in STD_LOGIC_VECTOR(1 downto 0);
	ETAJ_MINIM_MAXIM:in STD_LOGIC_VECTOR(3 downto 0);
	SENS_IN,CLOCK,SENZOR_USA,SENZOR_GREUTATE:in STD_LOGIC;
	ENABLE_DELETE,ENABLE_NUMARATOR_OUT:out STD_LOGIC;
	ETAJ_CURENT_OUT:out STD_LOGIC_VECTOR(3 downto 0));	
end entity AUTOMAT;


architecture F_AUTOMAT of AUTOMAT is

signal ENABLE_NUMARATOR_ETAJ,CLOCK_DIVIZAT:STD_LOGIC;
signal ETAJ_CURENT:STD_LOGIC_VECTOR(3 downto 0);


begin
	A1:entity work.NUMARATOR_ETAJ(F_NUMARATOR_ETAJ) PORT MAP (SENS_IN,ENABLE_NUMARATOR_ETAJ,CLOCK_DIVIZAT,ETAJ_CURENT);															   
	A2:entity work.OPRIRE(F_OPRIRE) PORT MAP (ETAJ_CURENT,ETAJ_MINIM_MAXIM,INFORMATIE_IN,SENS_IN,CLOCK,SENZOR_USA,SENZOR_GREUTATE,ENABLE_NUMARATOR_ETAJ,ENABLE_DELETE);
	A3:entity work.DIVIZOR_1_SEC(F_DIVIZOR_1_SEC) PORT MAP (CLOCK,CLOCK_DIVIZAT);	
	ETAJ_CURENT_OUT <= ETAJ_CURENT;
	ENABLE_NUMARATOR_OUT <= ENABLE_NUMARATOR_ETAJ;
	
end architecture F_AUTOMAT;

