library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.STD_LOGIC_UNSIGNED.all;
--use IEEE.STD_LOGIC_ARITH.all;
use ieee.numeric_std.all;

entity TOP is
	port(ETAJ:in STD_LOGIC_VECTOR(3 downto 0);
	SUS,JOS,INTERIOR,SENZOR_GREUTATE,SENZOR_USA,CLOCK:in STD_LOGIC;
	USI_DESCHISE:out STD_LOGIC;
	INFORMATIE_OUT,INFORMATIE_INPUT:out STD_LOGIC_VECTOR(1 downto 0);
	ANOD,ETAJ_MINIM_MAXIM_OUT:out STD_LOGIC_VECTOR(3 downto 0);
	CATOD:out STD_LOGIC_VECTOR(6 downto 0));
end entity TOP;


architecture F_TOP of TOP is

signal WE,SENS,ENABLE_DELETE,ENABLE_NUMARATOR,CLOCK_DIVIZAT:STD_LOGIC;
signal INFORMATIE_AUTOMAT,INFORMATIE_MEMORIE:STD_LOGIC_VECTOR(1 downto 0);
signal ETAJ_MINIM_MAXIM,ETAJ_CURENT,ETAJ_ADAUGARE:STD_LOGIC_VECTOR(3 downto 0);


begin
	T1:entity work.AUTOMAT(F_AUTOMAT) PORT MAP (INFORMATIE_AUTOMAT,ETAJ_MINIM_MAXIM,SENS,CLOCK,SENZOR_USA,SENZOR_GREUTATE,ENABLE_DELETE,ENABLE_NUMARATOR,ETAJ_CURENT);
	T2:entity work.INPUT(F_INPUT) PORT MAP (ETAJ,ETAJ_CURENT,SUS,JOS,INTERIOR,WE,ETAJ_ADAUGARE,INFORMATIE_MEMORIE);
	T3:entity work.MEMORIE(F_MEMORIE) PORT MAP (WE,ENABLE_DELETE,CLOCK_DIVIZAT,ETAJ_ADAUGARE,ETAJ_CURENT,INFORMATIE_MEMORIE,INFORMATIE_AUTOMAT,ETAJ_MINIM_MAXIM,SENS);
	T4:entity work.AFISARE(F_AFISARE) PORT MAP (ETAJ_CURENT,CLOCK,CATOD,ANOD);
	T5:entity work.DIVIZOR_1_SEC(F_DIVIZOR_1_SEC) PORT MAP (CLOCK,CLOCK_DIVIZAT);
	
	
	INFORMATIE_INPUT <= INFORMATIE_MEMORIE;
	INFORMATIE_OUT <= INFORMATIE_AUTOMAT;
	ETAJ_MINIM_MAXIM_OUT <= ETAJ_MINIM_MAXIM;
	USI_DESCHISE <= not(ENABLE_NUMARATOR);	
end architecture F_TOP;